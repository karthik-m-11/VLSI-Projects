// pkg/defines.svh
`ifndef DEFINES_SVH
`define DEFINES_SVH

// APB parameters
`define ADDR_WIDTH 16
`define DATA_WIDTH 32
`define MEM_DEPTH  256

// Verbosity levels
`define VERBOSITY UVM_MEDIUM

// Error codes
`define ERR_INVALID_ADDR 1

`endif